`include "frameSequencer.v"

module frameSequencerTest();


endmodule
